module num

pub fn add(x int, y int) int {
    return x + y
}